module font_rom ( input [9:0]	addr,
						output [63:0]	data
					 );

	parameter ADDR_WIDTH = 10;
   parameter DATA_WIDTH =  64;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	
         // code x00
        64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, // 0	  
        64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  // 1	  
        64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  // 2		  
        64'b0000000011111111111111110000000011111111111111110000000000000000, 
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,    
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000, // 3 		  
		  64'b0000000011111111111111110000000011111111111111110000000000000000, 
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,    
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000, // 4	  
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000, //5		  
		  64'b0000000011111111111111110000000011111111111111110000000000000000, 
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,    
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000, // 6		  
		  64'b0000000011111111111111110000000011111111111111110000000000000000, 
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,    
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000, // 7
		  64'b0000000011111111111111110000000011111111111111110000000000000000, 
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,    
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000, // 8
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000, //9
		  64'b0000000011111111111111110000000011111111111111110000000000000000, 
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,    
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000, // 10
		  64'b0000000011111111111111110000000011111111111111110000000000000000, 
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,    
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000, // 11
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, // 12
        64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  // 13
        64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  // 14 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  // 15
         //A code x01
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
        64'b0000000000000000000000001111111100000000000000000000000000000000,
		  64'b0000000000000000000000001111111100000000000000000000000000000000,
		  64'b0000000000000000000000001111111100000000000000000000000000000000,
		  64'b0000000000000000000000001111111100000000000000000000000000000000,
		  64'b0000000000000000000000001111111100000000000000000000000000000000,
		  64'b0000000000000000000000001111111100000000000000000000000000000000,
		  64'b0000000000000000000000001111111100000000000000000000000000000000,
		  64'b0000000000000000000000001111111100000000000000000000000000000000,
        64'b0000000000000000111111111111111111111111000000000000000000000000,
		  64'b0000000000000000111111111111111111111111000000000000000000000000,
		  64'b0000000000000000111111111111111111111111000000000000000000000000,
		  64'b0000000000000000111111111111111111111111000000000000000000000000,
		  64'b0000000000000000111111111111111111111111000000000000000000000000,
		  64'b0000000000000000111111111111111111111111000000000000000000000000,
		  64'b0000000000000000111111111111111111111111000000000000000000000000,
		  64'b0000000000000000111111111111111111111111000000000000000000000000,
        64'b0000000011111111111111110000000011111111111111110000000000000000,
		  64'b0000000011111111111111110000000011111111111111110000000000000000,
		  64'b0000000011111111111111110000000011111111111111110000000000000000,
		  64'b0000000011111111111111110000000011111111111111110000000000000000,
		  64'b0000000011111111111111110000000011111111111111110000000000000000,
		  64'b0000000011111111111111110000000011111111111111110000000000000000,
		  64'b0000000011111111111111110000000011111111111111110000000000000000,
		  64'b0000000011111111111111110000000011111111111111110000000000000000,
		  64'b0000000011111111111111110000000011111111111111110000000000000000,
        64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
        64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
        64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
         // code x02
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //0
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //1  
		  64'b1111111111111111111111111111111111111111111111110000000000000000,
		  64'b1111111111111111111111111111111111111111111111110000000000000000,
		  64'b1111111111111111111111111111111111111111111111110000000000000000,
		  64'b1111111111111111111111111111111111111111111111110000000000000000,
		  64'b1111111111111111111111111111111111111111111111110000000000000000,
		  64'b1111111111111111111111111111111111111111111111110000000000000000,
		  64'b1111111111111111111111111111111111111111111111110000000000000000,
		  64'b1111111111111111111111111111111111111111111111110000000000000000, //2  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, 
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,    
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, // 3		  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, 
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,    
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, // 4
		  64'b0000000011111111111111110000000000000000111111111111111100000000, 
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,    
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, // 5
		  64'b0000000011111111111111111111111111111111111111110000000000000000, 
		  64'b0000000011111111111111111111111111111111111111110000000000000000,  
		  64'b0000000011111111111111111111111111111111111111110000000000000000,    
		  64'b0000000011111111111111111111111111111111111111110000000000000000,  
		  64'b0000000011111111111111111111111111111111111111110000000000000000,  
		  64'b0000000011111111111111111111111111111111111111110000000000000000,  
		  64'b0000000011111111111111111111111111111111111111110000000000000000,  
		  64'b0000000011111111111111111111111111111111111111110000000000000000, // 6
		  64'b0000000011111111111111110000000000000000111111111111111100000000, 
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,    
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, // 7
		  64'b0000000011111111111111110000000000000000111111111111111100000000, 
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,    
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, // 8
		  64'b0000000011111111111111110000000000000000111111111111111100000000, 
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,    
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, // 9
		  64'b0000000011111111111111110000000000000000111111111111111100000000, 
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,    
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, // a
		  64'b1111111111111111111111111111111111111111111111110000000000000000,
		  64'b1111111111111111111111111111111111111111111111110000000000000000,
		  64'b1111111111111111111111111111111111111111111111110000000000000000,
		  64'b1111111111111111111111111111111111111111111111110000000000000000,
		  64'b1111111111111111111111111111111111111111111111110000000000000000,
		  64'b1111111111111111111111111111111111111111111111110000000000000000,
		  64'b1111111111111111111111111111111111111111111111110000000000000000,
		  64'b1111111111111111111111111111111111111111111111110000000000000000, //b
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //d
        64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //e
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //f
        //C  x03
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
        64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
        64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
        64'b1111111111111111000000000000000000000000000000001111111100000000,
		  64'b1111111111111111000000000000000000000000000000001111111100000000,
		  64'b1111111111111111000000000000000000000000000000001111111100000000,
		  64'b1111111111111111000000000000000000000000000000001111111100000000,
		  64'b1111111111111111000000000000000000000000000000001111111100000000,
		  64'b1111111111111111000000000000000000000000000000001111111100000000,
		  64'b1111111111111111000000000000000000000000000000001111111100000000,
		  64'b1111111111111111000000000000000000000000000000001111111100000000,
        64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
        64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
        64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
         // code x04
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //0
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //1	
		  64'b1111111111111111111111111111111111111111000000000000000000000000,
		  64'b1111111111111111111111111111111111111111000000000000000000000000,
		  64'b1111111111111111111111111111111111111111000000000000000000000000,
		  64'b1111111111111111111111111111111111111111000000000000000000000000,
		  64'b1111111111111111111111111111111111111111000000000000000000000000,
		  64'b1111111111111111111111111111111111111111000000000000000000000000,
		  64'b1111111111111111111111111111111111111111000000000000000000000000,
		  64'b1111111111111111111111111111111111111111000000000000000000000000, //2 
		  64'b0000000011111111111111110000000011111111111111110000000000000000, 
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,    
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000, // 3
		  64'b0000000011111111111111110000000000000000111111111111111100000000, 
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,    
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, // 4
		  64'b0000000011111111111111110000000000000000111111111111111100000000, 
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,    
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, // 5
		  64'b0000000011111111111111110000000000000000111111111111111100000000, 
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,    
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, // 6
		  64'b0000000011111111111111110000000000000000111111111111111100000000, 
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,    
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, // 7
		  64'b0000000011111111111111110000000000000000111111111111111100000000, 
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,    
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, // 8
		  64'b0000000011111111111111110000000000000000111111111111111100000000, 
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,    
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, // 9
		  64'b0000000011111111111111110000000011111111111111110000000000000000, 
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,    
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000,  
		  64'b0000000011111111111111110000000011111111111111110000000000000000, // a
		  64'b1111111111111111111111111111111111111111000000000000000000000000,
		  64'b1111111111111111111111111111111111111111000000000000000000000000,
		  64'b1111111111111111111111111111111111111111000000000000000000000000,
		  64'b1111111111111111111111111111111111111111000000000000000000000000,
		  64'b1111111111111111111111111111111111111111000000000000000000000000,
		  64'b1111111111111111111111111111111111111111000000000000000000000000,
		  64'b1111111111111111111111111111111111111111000000000000000000000000,
		  64'b1111111111111111111111111111111111111111000000000000000000000000, //b
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //d
        64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //e
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //f
        //0x05
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
        64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
        64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
        64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
        64'b0000000011111111111111110000000011111111000000000000000000000000,
		  64'b0000000011111111111111110000000011111111000000000000000000000000,
		  64'b0000000011111111111111110000000011111111000000000000000000000000,
		  64'b0000000011111111111111110000000011111111000000000000000000000000,
		  64'b0000000011111111111111110000000011111111000000000000000000000000,
		  64'b0000000011111111111111110000000011111111000000000000000000000000,
		  64'b0000000011111111111111110000000011111111000000000000000000000000,
		  64'b0000000011111111111111110000000011111111000000000000000000000000,
        64'b0000000011111111111111111111111111111111000000000000000000000000,
		  64'b0000000011111111111111111111111111111111000000000000000000000000,
		  64'b0000000011111111111111111111111111111111000000000000000000000000,
		  64'b0000000011111111111111111111111111111111000000000000000000000000,
		  64'b0000000011111111111111111111111111111111000000000000000000000000,
		  64'b0000000011111111111111111111111111111111000000000000000000000000,
		  64'b0000000011111111111111111111111111111111000000000000000000000000,
		  64'b0000000011111111111111111111111111111111000000000000000000000000,
        64'b0000000011111111111111110000000011111111000000000000000000000000,
		  64'b0000000011111111111111110000000011111111000000000000000000000000,
		  64'b0000000011111111111111110000000011111111000000000000000000000000,
		  64'b0000000011111111111111110000000011111111000000000000000000000000,
		  64'b0000000011111111111111110000000011111111000000000000000000000000,
		  64'b0000000011111111111111110000000011111111000000000000000000000000,
		  64'b0000000011111111111111110000000011111111000000000000000000000000,
		  64'b0000000011111111111111110000000011111111000000000000000000000000,
        64'b0000000011111111111111110000000000000000000000000000000000000000,
		  64'b0000000011111111111111110000000000000000000000000000000000000000,
		  64'b0000000011111111111111110000000000000000000000000000000000000000,
		  64'b0000000011111111111111110000000000000000000000000000000000000000,
		  64'b0000000011111111111111110000000000000000000000000000000000000000,
		  64'b0000000011111111111111110000000000000000000000000000000000000000,
		  64'b0000000011111111111111110000000000000000000000000000000000000000,
		  64'b0000000011111111111111110000000000000000000000000000000000000000,
        64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
		  64'b0000000011111111111111110000000000000000000000001111111100000000,
        64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
         // code x06
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //0
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //1
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000,
		  64'b1111111111111111111111111111111111111111111111111111111100000000, //2
		  64'b0000000011111111111111110000000000000000111111111111111100000000, 
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,    
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000,  
		  64'b0000000011111111111111110000000000000000111111111111111100000000, // 3
		  64'b0000000011111111111111110000000000000000000000001111111100000000, 
		  64'b0000000011111111111111110000000000000000000000001111111100000000,  
		  64'b0000000011111111111111110000000000000000000000001111111100000000,    
		  64'b0000000011111111111111110000000000000000000000001111111100000000,  
		  64'b0000000011111111111111110000000000000000000000001111111100000000,  
		  64'b0000000011111111111111110000000000000000000000001111111100000000,  
		  64'b0000000011111111111111110000000000000000000000001111111100000000,  
		  64'b0000000011111111111111110000000000000000000000001111111100000000, // 4
		  64'b0000000011111111111111110000000011111111000000000000000000000000, 
		  64'b0000000011111111111111110000000011111111000000000000000000000000,  
		  64'b0000000011111111111111110000000011111111000000000000000000000000,    
		  64'b0000000011111111111111110000000011111111000000000000000000000000,  
		  64'b0000000011111111111111110000000011111111000000000000000000000000,  
		  64'b0000000011111111111111110000000011111111000000000000000000000000,  
		  64'b0000000011111111111111110000000011111111000000000000000000000000,  
		  64'b0000000011111111111111110000000011111111000000000000000000000000, // 5
		  64'b0000000011111111111111111111111111111111000000000000000000000000, 
		  64'b0000000011111111111111111111111111111111000000000000000000000000,  
		  64'b0000000011111111111111111111111111111111000000000000000000000000,    
		  64'b0000000011111111111111111111111111111111000000000000000000000000,  
		  64'b0000000011111111111111111111111111111111000000000000000000000000,  
		  64'b0000000011111111111111111111111111111111000000000000000000000000,  
		  64'b0000000011111111111111111111111111111111000000000000000000000000,  
		  64'b0000000011111111111111111111111111111111000000000000000000000000, // 6
		  64'b0000000011111111111111110000000011111111000000000000000000000000, 
		  64'b0000000011111111111111110000000011111111000000000000000000000000,  
		  64'b0000000011111111111111110000000011111111000000000000000000000000,    
		  64'b0000000011111111111111110000000011111111000000000000000000000000,  
		  64'b0000000011111111111111110000000011111111000000000000000000000000,  
		  64'b0000000011111111111111110000000011111111000000000000000000000000,  
		  64'b0000000011111111111111110000000011111111000000000000000000000000,  
		  64'b0000000011111111111111110000000011111111000000000000000000000000, // 7
		  64'b0000000011111111111111110000000000000000000000000000000000000000, 
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000,    
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000, // 8
		  64'b0000000011111111111111110000000000000000000000000000000000000000, 
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000,    
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000, // 9
		  64'b0000000011111111111111110000000000000000000000000000000000000000, 
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000,    
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000,  
		  64'b0000000011111111111111110000000000000000000000000000000000000000, // a
		  64'b1111111111111111111111111111111100000000000000000000000000000000, 
		  64'b1111111111111111111111111111111100000000000000000000000000000000,  
		  64'b1111111111111111111111111111111100000000000000000000000000000000,    
		  64'b1111111111111111111111111111111100000000000000000000000000000000,  
		  64'b1111111111111111111111111111111100000000000000000000000000000000,  
		  64'b1111111111111111111111111111111100000000000000000000000000000000,  
		  64'b1111111111111111111111111111111100000000000000000000000000000000,  
		  64'b1111111111111111111111111111111100000000000000000000000000000000, // b
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, // c
        64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //d
        64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //e
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000, 
		  64'b0000000000000000000000000000000000000000000000000000000000000000,  //f
        //0x07
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
        64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
		  64'b0000000000000000111111111111111111111111111111110000000000000000,
        64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
        64'b1111111111111111000000000000000000000000000000001111111100000000,
		  64'b1111111111111111000000000000000000000000000000001111111100000000,
		  64'b1111111111111111000000000000000000000000000000001111111100000000,
		  64'b1111111111111111000000000000000000000000000000001111111100000000,
		  64'b1111111111111111000000000000000000000000000000001111111100000000,
		  64'b1111111111111111000000000000000000000000000000001111111100000000,
		  64'b1111111111111111000000000000000000000000000000001111111100000000,
		  64'b1111111111111111000000000000000000000000000000001111111100000000,
        64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
		  64'b1111111111111111000000000000000000000000000000000000000000000000,
        64'b1111111111111111000000001111111111111111111111111111111100000000,
		  64'b1111111111111111000000001111111111111111111111111111111100000000,
		  64'b1111111111111111000000001111111111111111111111111111111100000000,
		  64'b1111111111111111000000001111111111111111111111111111111100000000,
		  64'b1111111111111111000000001111111111111111111111111111111100000000,
		  64'b1111111111111111000000001111111111111111111111111111111100000000,
		  64'b1111111111111111000000001111111111111111111111111111111100000000,
		  64'b1111111111111111000000001111111111111111111111111111111100000000,
        64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
		  64'b1111111111111111000000000000000000000000111111111111111100000000,
        64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
		  64'b0000000011111111111111110000000000000000111111111111111100000000,
        64'b0000000000000000111111111111111111111111000000001111111100000000,
		  64'b0000000000000000111111111111111111111111000000001111111100000000,
		  64'b0000000000000000111111111111111111111111000000001111111100000000,
		  64'b0000000000000000111111111111111111111111000000001111111100000000,
		  64'b0000000000000000111111111111111111111111000000001111111100000000,
		  64'b0000000000000000111111111111111111111111000000001111111100000000,
		  64'b0000000000000000111111111111111111111111000000001111111100000000,
		  64'b0000000000000000111111111111111111111111000000001111111100000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000,
		  64'b0000000000000000000000000000000000000000000000000000000000000000
		  
		  };


	assign data = ROM[addr];

endmodule  